module adder(a,b,result);
input[15:0] a,b;
output [15:0] result;
assign result = a+b;
endmodule